LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY GEN_ADD_SUB IS
    PORT ( DATA1_IN :  IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
           DATA2_IN :  IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
           RESULT   : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
           C        : OUT STD_LOGIC := '0'; 	-- CARR/BORROW
           OP       :  IN STD_LOGIC := '0'; 	-- 0 = ADD, 1 = SUB
           Z        : OUT STD_LOGIC := '0'; 	-- ZERO FLAG
           V        : OUT STD_LOGIC := '0');	-- OVERFLOW
END GEN_ADD_SUB;

ARCHITECTURE BEHAVIORAL OF GEN_ADD_SUB IS
  
  SIGNAL CARRYOUT : STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
  SIGNAL BUFF     : STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
  
BEGIN
 
 LSB : 
   ENTITY WORK.ADD_SUB(BEHAVIOR)
   PORT MAP(A => DATA1_IN(0), B => DATA2_IN(0), S => BUFF(0), CI => OP, CO => CARRYOUT(0));
   RESULT(0) <= BUFF(0);
 --   
 GEN : 
   FOR N IN 1 TO 30 GENERATE
     OTHER : ENTITY WORK.ADD_SUB(BEHAVIOR)
       PORT MAP(A => DATA1_IN(N), B => DATA2_IN(N), S => RESULT(N), CI => CARRYOUT(N - 1), 
               CO => CARRYOUT(N));
 END GENERATE GEN;
 --
 MSB : 
   ENTITY WORK.ADD_SUB(BEHAVIOR)
   PORT MAP(A => DATA1_IN(31), B => DATA2_IN(31), S => RESULT(31), CI => CARRYOUT(30), 
           CO => CARRYOUT(31)); 
 --		   
 C <= CARRYOUT(31);  
 V <= CARRYOUT(30) XOR CARRYOUT(31);
 Z <= '1' WHEN  BUFF = "00000000000000000000000000000000" ELSE '0';
END BEHAVIORAL;
