LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ALU IS
  PORT(Z            : OUT  STD_LOGIC := '0';
       O            : OUT  STD_LOGIC := '0';
       C            : OUT  STD_LOGIC := '0';
       EN           :  IN  STD_LOGIC := '0';
       ALUCTR       :  IN  STD_LOGIC_VECTOR(2  DOWNTO 0) := "000";
       RESULT_ALU   : OUT  STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
       READDATA1_ALU:  IN  STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
       READDATA2_ALU:  IN  STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000"
       );
END ALU;

ARCHITECTURE BEHAVIOR OF ALU IS
  
  SIGNAL DATA1 : STD_LOGIC_VECTOR(31 DOWNTO 0):= "00000000000000000000000000000000";
  SIGNAL DATA2 : STD_LOGIC_VECTOR(31 DOWNTO 0):= "00000000000000000000000000000000";
  
  BEGIN

    PROCESS(EN)
      BEGIN
        IF (EN = '1') THEN
          CASE ALUCTR IS
            WHEN "000" => -- ADDER
              READDATA1 <= R0;
            WHEN "001" => -- SUBBTRACTER
              READDATA1 <= R1;
            WHEN "010" => -- AND
              READDATA1 <= R2;
            WHEN "011" => -- OR
              READDATA1 <= R3;
            WHEN "100" => -- LOGIC SHIFT LEFT
              READDATA1 <= R4;
            WHEN "101" => -- LOGIC SHIFT RIGHT
              READDATA1 <= R5;
            WHEN "110" => -- ARITHMETIC SHIFT LEFT
              READDATA1 <= R6;
            WHEN "111" => -- ARITHMETIC SHIFT RIGHT
              READDATA1 <= R7;
            WHEN OTHERS =>
            END CASE;
      ELSE
        
      END IF; 
    END PROCESS;
    
	 
END BEHAVIOR;


