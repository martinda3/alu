LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 

ENTITY OPMUX_TB  IS 
END; 
 
ARCHITECTURE OPMUX_TB_ARCH OF OPMUX_TB IS

  SIGNAL SAL  :  STD_LOGIC := 'U'; 
  SIGNAL SLR  :  STD_LOGIC := 'U'; 
  SIGNAL ADD  :  STD_LOGIC := 'U'; 
  SIGNAL SAR  :  STD_LOGIC := 'U'; 
  SIGNAL SUB  :  STD_LOGIC := 'U'; 
  SIGNAL ORR  :  STD_LOGIC := 'U'; 
  SIGNAL ANDD :  STD_LOGIC := 'U'; 
  SIGNAL SLLL :  STD_LOGIC := 'U'; 
  SIGNAL OP   :  STD_LOGIC_VECTOR (2 DOWNTO 0) := "UUU"; 

  COMPONENT OPMUX  
    PORT ( 
      SAL  : OUT STD_LOGIC; 
      SLR  : OUT STD_LOGIC; 
      ADD  : OUT STD_LOGIC; 
      SAR  : OUT STD_LOGIC; 
      SUB  : OUT STD_LOGIC; 
      ORR  : OUT STD_LOGIC; 
      ANDD : OUT STD_LOGIC; 
      SLLL : OUT STD_LOGIC; 
      OP   : IN STD_LOGIC_VECTOR (2 DOWNTO 0)); 
  END COMPONENT ; 

BEGIN
  DUT  : OPMUX  
    PORT MAP ( 
      SAL  => SAL,
      SLR  => SLR,
      ADD  => ADD,
      SAR  => SAR,
      SUB  => SUB,
      ORR  => ORR,
      ANDD => ANDD,
      SLLL => SLLL,
      OP   => OP); 
END ; 

