LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY GEN_AND IS
    PORT ( DATA1_IN :  IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
           DATA2_IN :  IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
           RESULT   : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000");-- OVERFLOW
END GEN_AND;

ARCHITECTURE BEHAVIORAL OF GEN_AND IS
BEGIN      
 GEN : FOR N IN 0 TO 31 GENERATE
   OTHER : ENTITY WORK.BITAND(BEHAVIOR)
   PORT MAP(A => DATA1_IN(N), B => DATA2_IN(N), S => RESULT(N));
 END GENERATE GEN;
END BEHAVIORAL;
