library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity GEN_ADD_SUB is
    Port ( DATA1_IN :  in STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
           DATA2_IN :  in STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
           RESULT   : out STD_LOGIC_VECTOR(31 DOWNTO 0) := "UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU";
           C        : out STD_LOGIC := 'U'; -- CARR/BORROW
           OP       :  IN STD_LOGIC := '1'; -- 0 = ADD, 1 = SUB
           Z        : out STD_LOGIC := '0'; -- ZERO FLAG
           V        : out STD_LOGIC := 'U');-- OVERFLOW
end GEN_ADD_SUB;

architecture Behavioral of GEN_ADD_SUB is
  
  SIGNAL CARRYOUT : STD_LOGIC_VECTOR(32 DOWNTO 0) := "00000000000000000000000000000000U";
  SIGNAL BUFF     : STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
  SIGNAL Z_FLAG   : STD_LOGIC := '0';
  SIGNAL OUTPUT   : STD_LOGIC := 'U';
begin
 -- ADD OR SUB FLAG
 PROCESS(OP)
   BEGIN
 CARRYOUT(0) <= OP;
 END PROCESS;
 -- COMPONENT GENERATOR
 GEN : FOR N IN 31 DOWNTO 0 GENERATE
 -- ADDER SUBTRACTOR
 OTHER : ENTITY WORK.ADD_SUB(BEHAVIOR)
 PORT MAP(A => DATA1_IN(N), 
          B => DATA2_IN(N), 
          S => BUFF(N),      -- LOCAL SIGNAL TO UPDATE ZERO FLAG
          CI => CARRYOUT(N), 
          CO => CARRYOUT(N + 1));
 -- UPDATE ZERO FLAG
 Z_FLAG <= '1' WHEN OUTPUT = '1';
 END GENERATE GEN;
 -- FLAGS
 PROCESS(CARRYOUT(32))
   BEGIN
    RESULT(31 DOWNTO 0) <= BUFF(31 DOWNTO 0);
    C <= CARRYOUT(32);
    V <= CARRYOUT(32) XOR CARRYOUT(31);
    IF (Z_FLAG = '1') THEN
      Z <= '0';
   ELSE 
     Z <= '1';
   END IF;
 END PROCESS;
end Behavioral;
