LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY GEN_ARIGHT IS
    PORT ( DATA1_IN :  IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000100000000001";
           RESULT   : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000");
END GEN_ARIGHT;

ARCHITECTURE BEHAVIORAL OF GEN_ARIGHT IS

  SIGNAL HOLDER : STD_LOGIC_VECTOR(32 DOWNTO 0):= "000000000000000000000000000000000";
  
BEGIN  
    
 GEN : 
   FOR N IN 31 DOWNTO 1 GENERATE
   OTHER : 
     ENTITY WORK.SLEFT(BEHAVIOR)
     PORT MAP(A => DATA1_IN(N), S => HOLDER(N));
 END GENERATE GEN;
 --
 RESULT(30 DOWNTO 0) <= HOLDER(31 DOWNTO 1);
 RESULT(31) <= HOLDER(31);
END BEHAVIORAL;