LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL;
 
ENTITY ADDER_TB_ARCH IS 
END ADDER_TB_ARCH; 
 
ARCHITECTURE ADDER_TB_ARCH OF ADDER_TB IS 
  
  TYPE EN_ARRAY  IS ARRAY (1 TO 10) OF STD_LOGIC;
  TYPE REG_ARRAY IS ARRAY (1 TO 10) OF STD_LOGIC_VECTOR(2  DOWNTO 0);
  TYPE DATAARRAY IS ARRAY (1 TO 10) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
  
  CONSTANT DELAY    :  TIME := 10 NS;
  
  CONSTANT OP_IN    :  EN_ARRAY  := ('0',     '1',   '0',   '1',   '0',   '1',   '0',   '0',   '0',   '0');
  
  CONSTANT A_IN   :  DATAARRAY := ("00000000000000000000000000000000", "00000000000000000000000000000000",
                                    "00000000000000000000000000000000", "00000000000000000000000000000000",
                                    "11111111111111111111111111111111", "00000000000000000000000000000000",
                                    "00000000000000000000000000000000", "00000000000000000000000000000000",
                                    "00000000000000000000000000000000", "00000000000000000000000000000000");
                                     
  CONSTANT B_IN   :  DATAARRAY := ("00000000000000000000000000000000", "00000000000000000000000000000000",
                                     "00000000000000000000000000000000", "00000000000000000000000000000000",
                                     "00000000000000000000000000000000", "00000000000000000000000000000000",
                                     "00000000000000000000000000000000", "00000000000000000000000000000000",
                                     "00000000000000000000000000000000", "00000000000000000000000000000000");
  
  
  SIGNAL OP    :  STD_LOGIC := '0';
  SIGNAL COUT   :  STD_LOGIC := '0';
  SIGNAL SUM  :  STD_LOGIC_VECTOR (31 DOWNTO 0) := "00000000000000000000000000000000"; 
  SIGNAL A  :  STD_LOGIC_VECTOR (31 DOWNTO 0) := "00000000000000000000000000000000"; 
  SIGNAL B  :  STD_LOGIC_VECTOR (31 DOWNTO 0) := "00000000000000000000000000000000"; 
    
  COMPONENT REGISTER_FILE  
    PORT ( 
      OP   :  IN STD_LOGIC ; 
      COUT  :  IN STD_LOGIC ; 
      SUM :  IN STD_LOGIC_VECTOR (31 DOWNTO 0); 
      A : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      B : OUT STD_LOGIC_VECTOR (31 DOWNTO 0));  
  END COMPONENT; 
  
BEGIN   
 
  TEST : PROCESS
    VARIABLE I : INTEGER := 1;
    BEGIN
      FOR I IN 1 TO 10 LOOP
        OP   <= OP_IN(I);
        B <= B_IN(I);
        A <= A_IN(I);
        WAIT FOR DELAY;
      END LOOP;
      WAIT;
    END PROCESS TEST;
 
--  CHECK : PROCESS
--    VARIABLE I : INTEGER := 1;
--    BEGIN
--      FOR I IN 1 TO 10 LOOP
--        REGREAD   <= RR_IN(I);
--        REGWRITE  <= RW_IN(I);
--        REGS      <= RS_IN(I);
--        REGT      <= RT_IN(I);
--        REGD      <= RD_IN(I);
--        WRITEDATA <= WR_IN(I);
--        WAIT FOR DELAY/2;
--      END LOOP;
--      WAIT;
--    END PROCESS CHECK;

  DUT  : REGISTER_FILE  
    PORT MAP ( 
      REGREAD   => REGREAD,
      REGWRITE  => REGWRITE,
      REGS      => REGS,
      REGT      => REGT,
      REGD      => REGD,
      WRITEDATA => WRITEDATA,
      READDATA1 => READDATA1,
      READDATA2 => READDATA2) ; 
      
END ADDER_TB_ARCH; 

