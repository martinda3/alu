library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity GEN_ADD_SUB is
    Port ( DATA1_IN :  in STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000001";
           DATA2_IN :  in STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000001";
           RESULT   : out STD_LOGIC_VECTOR(31 DOWNTO 0) := "UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU";
           C        : out STD_LOGIC := 'U';
           OP       :  IN STD_LOGIC := '1';
           Z        : out STD_LOGIC := '0';
           V        : out STD_LOGIC := 'U');
end GEN_ADD_SUB;

architecture Behavioral of GEN_ADD_SUB is
  
  SIGNAL CARRYOUT : STD_LOGIC_VECTOR(32 DOWNTO 0) := "00000000000000000000000000000000U";
  SIGNAL Z_FLAG   : STD_LOGIC := '0';
  SIGNAL OUTPUT : STD_LOGIC := 'U';
begin
 CARRYOUT(0) <= OP;
 GEN : FOR N IN 31 DOWNTO 0 GENERATE
 OTHER : ENTITY WORK.ADD_SUB(BEHAVIOR)
 PORT MAP(A => DATA1_IN(N), B => DATA2_IN(N), S => OUTPUT, CI => CARRYOUT(N), CO => CARRYOUT(N + 1));
 RESULT(N) <= OUTPUT;
 Z_FLAG <= '1' WHEN OUTPUT = '1';
 END GENERATE GEN;
 C <= CARRYOUT(32);
 V <= CARRYOUT(32) XOR CARRYOUT(31);
 Z <= '0' when Z_FLAG = '1' else
      '1' when Z_FLAG = '0';
 
end Behavioral;
